package System_pkg;

import uvm_pkg::*;

`include "uvm_macros.svh"
`include "System_item.svh"
`include "System_sequencer.svh"
`include "System_driver.svh"
`include "System_monitor.svh"
`include "System_agent.svh"

    
endpackage: System_pkg