package APB_pkg;

import uvm_pkg::*;


`include "uvm_macros.svh"
`include "APB_item.svh"
`include "APB_driver.svh"
`include "APB_monitor.svh"
`include "APB_sequencer.svh"
`include "APB_agent.svh"
`include "Coverages_afvip.svh"



    
endpackage: APB_pkg