package Test_pkg;

import uvm_pkg::*;
import APB_pkg::*;
import System_pkg::*;
import AFVIP_pkg::*;

`include "uvm_macros.svh"
`include "APB_sequence.svh"
`include "System_sequence.svh"
`include "Test_scoreboard.svh"
`include "Test_enviroment.svh"
`include "afvip_test.svh"


    
endpackage: Test_pkg