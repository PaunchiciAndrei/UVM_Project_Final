package AFVIP_pkg;

import uvm_pkg::*;

`include "uvm_macros.svh"

`include "AFVIP_item.svh"
`include "AFVIP_monitor.svh"
`include "AFVIP_agent.svh"

endpackage: AFVIP_pkg